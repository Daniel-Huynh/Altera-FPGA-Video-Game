module Choose_Pattern(Clock, Reset, out);
	input logic Clock, Reset;
	output logic out;
			
endmodule